// $Id: $
// File name:   fir_filter.sv
// Created:     3/11/2021
// Author:      Ti-Wei Chen
// Lab Section: 337-06
// Version:     1.0  Initial Design Entry
// Description: Finite Impulse Response (FIR) Filter Design

module fir_filter
(
	input wire clk,
	input wire n_reset,
	input reg [15:0] sample_data,
	input reg [15:0] fir_coefficient,
	input reg load_coeff,
	input reg data_ready,
	output wire one_k_samples,
	output wire modwait,
	output wire [15:0] fir_out,
	output wire err
);

	reg sync_load_coeff;
	reg sync_data_ready;
	reg overflow;
	reg cnt_up;
	reg clear;
	reg [2:0] op;
	reg [3:0] src1;
	reg [3:0] src2;
	reg [3:0] dest;
	reg [16:0] outreg_data;

	sync_low SYNC_LR (.clk(clk), .n_rst(n_reset), .async_in(load_coeff), .sync_out(sync_load_coeff));

	sync_low SYNC_DR (.clk(clk), .n_rst(n_reset), .async_in(data_ready), .sync_out(sync_data_ready));

	counter COUNT (.clk(clk), .n_rst(n_reset), .cnt_up(cnt_up), .clear(clear), .one_k_samples(one_k_samples));

	controller CONTROL
	(
		.clk(clk),
		.n_rst(n_reset),
		.dr(sync_data_ready),
		.lc(sync_load_coeff),
		.overflow(overflow),
		.cnt_up(cnt_up),
		.clear(clear),
		.modwait(modwait),
		.op(op),
		.src1(src1),
		.src2(src2),
		.dest(dest),
		.err(err)
	);

	datapath DATAPATH
	(
		.clk(clk),
		.n_reset(n_reset),
		.op(op),
		.src1(src1),
		.src2(src2),
		.dest(dest),
		.ext_data1(sample_data),
		.ext_data2(fir_coefficient),
		.outreg_data(outreg_data),
		.overflow(overflow)
	);

	magnitude MAGNITUDE (.in(outreg_data), .out(fir_out));

endmodule
